(** Linear Scan Register Allocator

    The linear scan algorithm in this module is documented by the paper
    "Optimized Interval Splitting in a Linear Scan Register Allocator" by
    Christian Wimmer and Hanspeter Mӧssenbӧck:

    https://www.usenix.org/legacy/events/vee05/full_papers/p132-wimmer.pdf *)

Require Import Coq.Arith.EqNat.
Require Import Coq.Lists.List.
Require Import Coq.Numbers.Natural.Peano.NPeano.
Require Import Coq.Program.Basics.
Require Import Coq.Program.Tactics.
Require Import Coq.Logic.ProofIrrelevance.
Require Import Coq.Sorting.Sorting.
Require Import Coq.Structures.Orders.
Require Import Recdef.
Require Import Lib.
Require Import RState.
Require String.

Module Import LN := ListNotations.

Open Scope string_scope.
Open Scope nat_scope.
Open Scope program_scope.

Generalizable All Variables.

(****************************************************************************)

(** * Core data types *)

(** ** UsePos *)

(** A "use position", or [UsePos], identifies an exact point in the
    instruction stream where a particular variable is used.  If this usage
    requires the use of a physical register, then [regReq] is [true] for that
    use position. *)

Record UsePos : Set := {
  uloc   : nat;
  regReq : bool
}.

(** ** Range *)

(** The extent of a [Range] is the set of locations it ranges over.  By
    summing the extent of a list of ranges, we have an idea of how much ground
    is left to cover, and this gives us a notion of well-founded recursion for
    iterating over intervals that may split as we examine them -- i.e., whose
    total extent must decrease after each pass.

    A Range is built up from a set of use positions, and defines the inclusive
    range of those positions.  It can be extended, or split, but never shrunk.
    Also, the non-empty list of use positions is not guaranteed to be in any
    order, and overlapping use positions are accepted but only the most recent
    one "wins". *)

Record RangeDesc := {
    rbeg : nat;
    rend : nat;
    ups  : NonEmpty UsePos;

    range_nonempty : rbeg < rend         (* this comes in handy *)
}.

Inductive Range : RangeDesc -> Set :=
  | R_Sing u :
      Range {| rbeg := uloc u
             ; rend := S (uloc u)
             ; ups  := NE_Sing u
             ; range_nonempty := le_n (S (uloc u))
             |}
  | R_Cons u x : Range x -> forall (H : uloc u < rbeg x),
      Range {| rbeg := uloc u
             ; rend := rend x
             ; ups  := NE_Cons u (ups x)
             ; range_nonempty := Lt.lt_trans _ _ _ H (range_nonempty x)
             |}
  | R_Extend x b' e' : Range x ->
      Range {| rbeg := min b' (rbeg x)
             ; rend := Peano.max e' (rend x)
             ; ups  := ups x
             ; range_nonempty := min_lt_max _ _ _ _ (range_nonempty x)
             |}.

Definition rangeExtent (x : RangeDesc) := rend x - rbeg x.

Definition rangesIntersect `(x : RangeDesc) `(y : RangeDesc) : bool :=
  if rbeg x <? rbeg y
  then rbeg y <? rend x
  else rbeg x <? rend y.

Definition anyRangeIntersects (is js : NonEmpty RangeDesc) : bool :=
  fold_right
    (fun r b => orb b (existsb (rangesIntersect r) (NE_to_list js)))
    false (NE_to_list is).

(** ** Interval *)

(** A lifetime interval defines the lifetime of a variable.  It is defined as
    a list of ranges "covered" by that variable in the low-level intermediate
    representation (LIR).  Gaps in the list of ranges are called "lifetime
    holes".

    A lifetime is not necessarily only the distance that a variable is first
    and last used.  The lifetime of a variable used in a loop extends to the
    whole loop, for example, even if it is only used at the very end.  In this
    sense, coverage takes into account code flow, or what ranges would map to
    if all loops were unrolled, and then rolled back keeping track of
    coverage.

    Use positions are actual instructions where a variable is read from or
    written to, and whether it is required to be in a register at that
    point. *)

(** If for some reason we cannot assign a single register for all ranges, then
    the interval is split into two or more intervals, so each interval can be
    assigned its own register. *)

Record IntervalDesc := {
    ibeg : nat;
    iend : nat;
    rds  : NonEmpty RangeDesc;

    interval_nonempty : ibeg < iend         (* comes in handy *)
}.

Inductive Interval : IntervalDesc -> Set :=
  | I_Sing : forall x, Range x ->
      Interval {| ibeg := rbeg x
                ; iend := rend x
                ; rds  := NE_Sing x
                ; interval_nonempty := range_nonempty x
                |}
  | I_Cons1 : forall x y ib ie ne,
      Interval {| ibeg := ib; iend := ie; rds := NE_Sing y;
                  interval_nonempty := ne |}
        -> Range x -> forall (H : rend x <= ib),
      Interval {| ibeg := rbeg x
                ; iend := ie
                ; rds  := NE_Cons x (NE_Sing y)
                ; interval_nonempty := lt_le_shuffle (range_nonempty x) H ne
                |}
  | I_Consn : forall x y xs ib ie ne,
      Interval {| ibeg := ib; iend := ie; rds := NE_Cons y xs;
                  interval_nonempty := ne |}
        -> Range x -> forall (H : rend x <= ib),
      Interval {| ibeg := rbeg x
                ; iend := ie
                ; rds  := NE_Cons x (NE_Cons y xs)
                ; interval_nonempty := lt_le_shuffle (range_nonempty x) H ne
                |}.

Definition intervalStart `(i : Interval d) : nat := ibeg d.
Definition intervalEnd   `(i : Interval d) : nat := iend d.

Lemma Interval_nonempty : forall `(i : Interval rs),
  intervalStart i < intervalEnd i.
Proof.
  intros. unfold intervalStart, intervalEnd.
  induction i; simpl in *;
  induction r; simpl in *; min_max.
Qed.

Definition intervalCoversPos `(i : Interval rs) (pos : nat) : bool :=
  andb (intervalStart i <=? pos) (pos <? intervalEnd i).

Definition intervalExtent `(i : Interval rs) :=
  intervalEnd i - intervalStart i.

Lemma Interval_extent_nonempty : forall `(i : Interval rs),
  intervalExtent i > 0.
Proof.
  intros.
  unfold intervalExtent.
  pose (Interval_nonempty i).
  apply lt_minus in l. assumption.
Qed.

(****************************************************************************)

(** * Main algorithm *)

Section Allocator.

Variable maxReg : nat.          (* max number of registers *)

Hypothesis registers_exist : maxReg > 0.

Definition VirtReg := nat.
Definition PhysReg := fin maxReg.

(** ** ScanState *)

(** A [ScanState] is always relative to a current position (pos) as we move
    through the sequentialized instruction stream over which registers are
    allocated.. *)

Record ScanStateDesc := {
    nextInterval : nat;
    IntervalId   := fin nextInterval;

    unhandledExtent : nat;

    unhandled : list IntervalId;   (* starts after pos *)
    active    : list IntervalId;   (* ranges over pos *)
    inactive  : list IntervalId;   (* falls in lifetime hole *)
    handled   : list IntervalId;   (* ends before pos *)

    getInterval  : IntervalId -> { d : IntervalDesc & Interval d };
    assignments  : IntervalId -> option PhysReg;

    unhandled_sorted : LocallySorted cmp_le unhandled;

    all_state_lists  := unhandled ++ active ++ inactive ++ handled;
    lists_are_unique : NoDup all_state_lists
}.

Definition transportId `(H : nextInterval st <= nextInterval st')
  (x : IntervalId st) : IntervalId st'.
Proof.
  destruct st. destruct st'.
  unfold IntervalId0, IntervalId1 in *.
  unfold IntervalId in *. simpl in *.
  apply (fin_transport nextInterval0 nextInterval1 H).
  assumption.
Defined.

Lemma NoDup_wip : forall n x unh act inact hnd,
  NoDup (unh ++ act ++ inact ++ hnd) ->
  NoDup ((x :: map (fin_bump n) unh) ++
         map (fin_bump n) act ++ map (fin_bump n) inact ++
         map (fin_bump n) hnd).
Proof.
Admitted.

Lemma LocallySorted_fin_bump : forall n (x : fin (S n)) (xs : list (fin n)),
  LocallySorted cmp_le xs
    -> x = ultimate_Sn n
    -> LocallySorted cmp_le (x :: map (fin_bump n) xs).
Proof.
Admitted.

Lemma move_active_to_inactive : forall sd x,
  NoDup (unhandled sd ++ active sd ++ inactive sd ++ handled sd)
    -> In x (active sd)
    -> NoDup (unhandled sd ++ remove cmp_eq_dec x (active sd) ++
              (x :: inactive sd) ++ handled sd).
Proof.
  intros.
  apply NoDup_swap.
  rewrite <- app_assoc.
  rewrite <- app_assoc.
  apply NoDup_juggle.
  rewrite app_assoc.
  rewrite app_assoc.
  apply NoDup_swap.
  rewrite <- app_assoc.
  assumption.
  apply H0.
Defined.

Lemma move_active_to_handled : forall sd x,
  NoDup (unhandled sd ++ active sd ++ inactive sd ++ handled sd)
    -> In x (active sd)
    -> NoDup (unhandled sd ++ remove cmp_eq_dec x (active sd) ++
              inactive sd ++ x :: handled sd).
Proof.
  intros.
  apply NoDup_swap.
  rewrite <- app_assoc.
  rewrite <- app_assoc.
  apply NoDup_swap2.
  rewrite <- app_assoc.
  apply NoDup_juggle.
  rewrite app_assoc.
  apply NoDup_swap2.
  rewrite app_assoc.
  apply NoDup_swap.
  rewrite <- app_assoc.
  rewrite app_assoc.
  apply NoDup_swap2.
  rewrite <- app_assoc.
  assumption.
  apply H0.
Defined.

Definition move_inactive_to_active : forall sd x,
  NoDup (unhandled sd ++ active sd ++ inactive sd ++ handled sd)
    -> In x (inactive sd)
    -> NoDup (unhandled sd ++ x :: active sd ++
              remove cmp_eq_dec x (inactive sd) ++ handled sd).
Proof.
Admitted.

Definition move_inactive_to_handled : forall sd x,
  NoDup (unhandled sd ++ active sd ++ inactive sd ++ handled sd)
    -> In x (inactive sd)
    -> NoDup (unhandled sd ++ active sd ++
              remove cmp_eq_dec x (inactive sd) ++ x :: handled sd).
Proof.
Admitted.

(** The [ScanState] inductive data type describes the allowable state
    transitions that can be applied to a [ScanStateDesc] value.

    In essence there are five mutating operations:

    1. Create a new unhandled interval.  This can occur for two reasons:

       a. Adding a new interval to be considered before the linear scan
          algorithm has started.
       b. Splitting the current interval, which pushes back its "pieces" as
          new unhandled intervals.

    2. Remove the first unhandled interval.  This happens when we remove it in
       order to make it the new current interval.

    3. Add the current interval to the active list.

    4. Move an item from the active list to the inactive or handled lists.

    5. Move an item from the inactive list to the active or handled lists. *)

Inductive ScanState : ScanStateDesc -> Set :=
  | ScanState_nil :
    ScanState
      {| nextInterval     := 0
       ; unhandledExtent  := 0
       ; unhandled        := nil
       ; active           := nil
       ; inactive         := nil
       ; handled          := nil
       ; getInterval      := fin_contra
       ; assignments      := fin_contra
       ; unhandled_sorted := LSorted_nil _
       ; lists_are_unique := NoDup_nil _
       |}

  | ScanState_newUnhandled
      ni ue unh unhsort act inact hnd geti assgn lau :
    forall `(i : Interval d),
    ScanState
      {| nextInterval     := ni
       ; unhandledExtent  := ue
       ; unhandled        := unh
       ; active           := act
       ; inactive         := inact
       ; handled          := hnd
       ; getInterval      := geti
       ; assignments      := assgn
       ; unhandled_sorted := unhsort
       ; lists_are_unique := lau
       |} ->
    forall newi (H : newi = ultimate_Sn ni),
    ScanState
      {| nextInterval     := S ni
       ; unhandledExtent  := ue + intervalExtent i
       ; unhandled        := newi :: map (fin_bump ni) unh
       ; active           := map (fin_bump ni) act
       ; inactive         := map (fin_bump ni) inact
       ; handled          := map (fin_bump ni) hnd
       ; getInterval      :=
         fun n => match cmp_eq_dec n newi with
                  | left _ => existT _ d i
                  | right Hn => geti (fin_safe_reduce n (rew_in_not_eq H Hn))
                  end
       ; assignments      :=
         fun n => match cmp_eq_dec n newi with
                  | left _ => None
                  | right Hn => assgn (fin_safe_reduce n (rew_in_not_eq H Hn))
                  end
       ; unhandled_sorted := LocallySorted_fin_bump _ _ _ unhsort H
       ; lists_are_unique := NoDup_wip ni newi unh _ _ _ lau
       |}

  | ScanState_dropUnhandled
      ni ue x unh unhsort act inact hnd geti assgn lau :
    ScanState
      {| nextInterval     := ni
       ; unhandledExtent  := intervalExtent (projT2 (geti x)) + ue
       ; unhandled        := x :: unh
       ; active           := act
       ; inactive         := inact
       ; handled          := hnd
       ; getInterval      := geti
       ; assignments      := assgn
       ; unhandled_sorted := unhsort
       ; lists_are_unique := lau
       |} ->
    ScanState
      {| nextInterval     := ni
       ; unhandledExtent  := ue
       ; unhandled        := unh
       ; active           := act
       ; inactive         := inact
       ; handled          := hnd
       ; getInterval      := geti
       ; assignments      := assgn
       ; unhandled_sorted := LocallySorted_uncons _ _ _ _ unhsort
       ; lists_are_unique := NoDup_uncons _ _ _ _ lau
       |}

  | ScanState_moveActiveToInactive sd x :
    ScanState sd -> forall (H : In x (active sd)),
    ScanState
      {| nextInterval     := nextInterval sd
       ; unhandledExtent  := unhandledExtent sd
       ; unhandled        := unhandled sd
       ; active           := remove cmp_eq_dec x (active sd)
       ; inactive         := x :: inactive sd
       ; handled          := handled sd
       ; getInterval      := getInterval sd
       ; assignments      := assignments sd
       ; unhandled_sorted := unhandled_sorted sd
       ; lists_are_unique := move_active_to_inactive sd x (lists_are_unique sd) H
       |}

  | ScanState_moveActiveToHandled sd x :
    ScanState sd -> forall (H : In x (active sd)),
    ScanState
      {| nextInterval     := nextInterval sd
       ; unhandledExtent  := unhandledExtent sd
       ; unhandled        := unhandled sd
       ; active           := remove cmp_eq_dec x (active sd)
       ; inactive         := inactive sd
       ; handled          := x :: handled sd
       ; getInterval      := getInterval sd
       ; assignments      := assignments sd
       ; unhandled_sorted := unhandled_sorted sd
       ; lists_are_unique := move_active_to_handled sd x (lists_are_unique sd) H
       |}

  | ScanState_moveInactiveToActive sd x :
    ScanState sd -> forall (H : In x (inactive sd)),
    ScanState
      {| nextInterval     := nextInterval sd
       ; unhandledExtent  := unhandledExtent sd
       ; unhandled        := unhandled sd
       ; active           := x :: active sd
       ; inactive         := remove cmp_eq_dec x (inactive sd)
       ; handled          := handled sd
       ; getInterval      := getInterval sd
       ; assignments      := assignments sd
       ; unhandled_sorted := unhandled_sorted sd
       ; lists_are_unique := move_inactive_to_active sd x (lists_are_unique sd) H
       |}

  | ScanState_moveInactiveToHandled sd x :
    ScanState sd -> forall (H : In x (inactive sd)),
    ScanState
      {| nextInterval     := nextInterval sd
       ; unhandledExtent  := unhandledExtent sd
       ; unhandled        := unhandled sd
       ; active           := active sd
       ; inactive         := remove cmp_eq_dec x (inactive sd)
       ; handled          := x :: handled sd
       ; getInterval      := getInterval sd
       ; assignments      := assignments sd
       ; unhandled_sorted := unhandled_sorted sd
       ; lists_are_unique := move_inactive_to_handled sd x (lists_are_unique sd) H
       |}.

Tactic Notation "ScanState_cases" tactic(first) ident(c) :=
  first;
  [ Case_aux c "ScanState_nil"
  | Case_aux c "ScanState_newUnhandled"
  | Case_aux c "ScanState_dropUnhandled"
  | Case_aux c "ScanState_moveActiveToInactive"
  | Case_aux c "ScanState_moveActiveToHandled"
  | Case_aux c "ScanState_moveInactiveToActive"
  | Case_aux c "ScanState_moveInactiveToHandled"
  ].

Theorem ScanState_active_bounded : forall st,
  length (active st) <= nextInterval st.
Proof.
  destruct st. simpl.
  unfold all_state_lists0 in lists_are_unique0.
  compute.
  apply NoDup_unapp in lists_are_unique0.
  inversion lists_are_unique0.
  apply NoDup_swap in H0.
  apply NoDup_unapp in H0.
  inversion H0.
  apply fin_list in H2.
  auto.
Qed.

Ltac cmp_reflexive :=
  match goal with
    [ |- context [match cmp_eq_dec ?X ?X with _ => _ end] ] =>
      assert (cmp_eq_dec X X = left eq_refl) as Hrcmp
        by (intros; destruct (cmp_eq_dec X X);
              [ f_equal; apply proof_irrelevance
              | intuition ]);
      rewrite Hrcmp in *; clear Hrcmp; simpl in *
  end.

Theorem ScanState_unhandledExtent `(st : ScanState sd) :
  let unh := unhandled sd in
  let ue := unhandledExtent sd in
  IF unh = []
  then ue = 0
  else (forall i,
        let ie := intervalExtent (projT2 (getInterval sd i)) in
        IF unh = [i] then ue = ie else ue > ie).
Proof.
  ScanState_cases (induction st) Case; simpl in *.
  - Case "ScanState_nil". left. auto.
  - Case "ScanState_newUnhandled".
    right. split.
      apply not_eq_sym.
      apply nil_cons.
    intros. intuition.
    destruct unh eqn:Heqe; simpl.
      destruct (@cmp_eq_dec (fin (S ni)) (@fin_CompareSpec (S ni))
                            i0 newi) eqn:Heqe2.
        left. split. rewrite e. reflexivity.
        inversion IHst; inversion H0.
          simpl. omega.
        contradiction H1. reflexivity.
      admit.
    right. split.
      intuition. inversion H0.
    destruct (@cmp_eq_dec (fin (S ni)) (@fin_CompareSpec (S ni))
                          i0 newi) eqn:Heqe2.
      inversion IHst; inversion H0. inversion H1.
      simpl in *.
      specialize (H2 i0).
      contradiction H1. reflexivity.
    
    inversion IHst.
      destruct unh eqn:Heqe; simpl.
        right. split.
          unfold not. intros.
          inversion H1.
        intros.
        destruct (@cmp_eq_dec (fin (S ni)) (@fin_CompareSpec (S ni))
                              i0 newi) eqn:Heqe2.
          left. split. rewrite e. reflexivity.
          inversion H0. simpl. omega.
        right. split.
          unfold not in *. intros.
          apply n. congruence.
        
    destruct unh eqn:Heqe; simpl.
      right. split.
        unfold not. intros. inversion H0.
      intros. simpl in *.
      right. split.
        unfold not in *. intros.
        apply n. congruence.
      inversion IHst; inversion H0.
        rewrite H2 in *. simpl in *.
      rewrite Heqe2.
    admit.
  - Case "ScanState_dropUnhandled". admit.
  - Case "ScanState_moveActiveToInactive". admit.
  - Case "ScanState_moveActiveToHandled". admit.
  - Case "ScanState_moveInactiveToActive". admit.
  - Case "ScanState_moveInactiveToHandled". admit.
Admitted.

(** ** SSMorph *)

(** A [SSMorph] is a relation describe a lawful transition between two
    states.  It is a [PreOrder] relation. *)

Record SSMorph (sd1 : ScanStateDesc) (sd2 : ScanStateDesc) := {
    next_interval_increases : nextInterval sd1     <= nextInterval sd2;
    total_extent_decreases  : unhandledExtent sd2  <= unhandledExtent sd1;
    handled_count_increases : length (handled sd1) <= length (handled sd2)
}.

Arguments next_interval_increases [sd1 sd2] _.
Arguments total_extent_decreases  [sd1 sd2] _.
Arguments handled_count_increases [sd1 sd2] _.

Definition newSSMorph (s : ScanStateDesc) : SSMorph s s.
Proof. constructor; auto. Defined.

Program Instance SSMorph_PO : PreOrder SSMorph.
Obligation 1. constructor; auto. Defined.
Obligation 2.
  constructor; destruct H; destruct H0.
  transitivity (nextInterval y); auto.
  transitivity (unhandledExtent y); auto.
  transitivity (length (handled y)); auto.
Defined.

(** ** CurrentInterval *)

Record CurrentInterval `(st : ScanState sd) := {
    currentIntervalId : IntervalId sd;
    currentDesc       : IntervalDesc;
    currentInterval   : Interval currentDesc

    (* not_present : ~ In currentIntervalId (all_state_lists sd) *)
}.

Arguments currentIntervalId [sd st] _.
Arguments currentDesc       [sd st] _.
Arguments currentInterval   [sd st] _.

Record SSMorphSt (sd1 : ScanStateDesc) (sd2 : ScanStateDesc) : Prop := {
    is_SSMorph :> SSMorph sd1 sd2;

    total_extent_measurably_decreases :
      unhandledExtent sd2 < unhandledExtent sd1
}.

Program Instance SSMorphSt_Trans : Transitive SSMorphSt.
Obligation 1.
  constructor.
    destruct H. destruct H0.
    transitivity y; assumption.
  inversion H. inversion H0.
  destruct total_extent_measurably_decreases1. omega.
  destruct total_extent_measurably_decreases0. omega.
  right. omega.
Qed.

Theorem compose_SSMorph_with_SSMorphSt : forall (sd1 sd2 sd3 : ScanStateDesc),
  SSMorphSt sd1 sd2 -> SSMorph sd2 sd3 -> SSMorphSt sd1 sd3.
Proof.
  intros.
  constructor.
  inversion H.
  transitivity sd2; assumption.
  inversion H. inversion H0. omega.
Qed.

Theorem SSMorphSt_proj_unhandledExtent : forall (sd1 sd3 : ScanStateDesc),
  SSMorphSt sd1 sd3 -> unhandledExtent sd3 < unhandledExtent sd1.
Proof. intros. inversion H. assumption. Qed.

Lemma ScanState_unhandledExtent_nonzero `(st : ScanState sd) :
  length (unhandled sd) > 0 <-> unhandledExtent sd > 0.
Proof.
  intros.
  ScanState_cases (induction st) Case; simpl in *.
  - Case "ScanState_nil".
    split; intros; inversion H.
  - Case "ScanState_newUnhandled".
    pose (Interval_extent_nonempty i); omega.
  - Case "ScanState_dropUnhandled".
    apply ScanState_unhandledExtent in st.
    rename st into i. simpl in *.
    destruct unh eqn:Heqe.
      split; intros. inversion H.
      inversion i; inversion H0.
        inversion H1.
      specialize (H2 x).
      inversion H2; inversion H3.
        apply plus_eq_zero in H5. omega.
      contradiction H4. reflexivity.
    inversion i; inversion H.
      inversion H0.
    specialize (H1 x).
    inversion H1; inversion H2.
      split; intros; inversion H3.
    split; intros.
      apply plus_gt_zero in H4.
      assumption.
    simpl. apply Gt.gt_Sn_O.
  - Case "ScanState_moveActiveToInactive".  apply IHst.
  - Case "ScanState_moveActiveToHandled".   apply IHst.
  - Case "ScanState_moveInactiveToActive".  apply IHst.
  - Case "ScanState_moveInactiveToHandled". apply IHst.
Qed.

Lemma ScanState_no_unhandledExtent `(st : ScanState sd)
  (H : length (unhandled sd) = 0) : unhandledExtent sd = 0.
Proof.
  ScanState_cases (induction st) Case; simpl in *.
  - Case "ScanState_nil". apply H.
  - Case "ScanState_newUnhandled". inversion H.
  - Case "ScanState_dropUnhandled".
    apply ScanState_unhandledExtent in st.
    rename st into Hi. simpl in *.
    destruct unh eqn:Heqe.
      subst. inversion Hi; inversion H0. omega.
      apply nil_list_0 in H.
      specialize (H2 x).
      inversion H2; inversion H3. omega.
      contradiction H4. reflexivity.
    inversion H.
  - Case "ScanState_moveActiveToInactive".  apply IHst. assumption.
  - Case "ScanState_moveActiveToHandled".   apply IHst. assumption.
  - Case "ScanState_moveInactiveToActive".  apply IHst. assumption.
  - Case "ScanState_moveInactiveToHandled". apply IHst. assumption.
Defined.

Lemma ScanState_sole_unhandledExtent `(st : ScanState sd)
  (H : length (unhandled sd) = 1) :
  intervalExtent (projT2 (getInterval sd
                  (safe_hd (unhandled sd) (one_gt_zero _ H)))) =
  unhandledExtent sd.
Proof.
  pose proof st as Hi.
  apply ScanState_unhandledExtent in Hi.
  ScanState_cases (induction st) Case; simpl in *.
  - Case "ScanState_nil". inversion H.
  - Case "ScanState_newUnhandled".
    clear IHst.
    cmp_reflexive.
    inversion H.
    rewrite map_length in H2.
    pose (ScanState_no_unhandledExtent st). simpl in e.
    rewrite e; auto.
  - Case "ScanState_dropUnhandled".
    clear IHst.
    destruct unh eqn:Heqe. inversion H.
    assert (l = []). apply nil_list_0. auto.
    simpl in *. subst.
    inversion Hi; inversion H0. inversion H1.
    specialize (H2 f).
    inversion H2; inversion H3. auto.
    contradiction H4. reflexivity.
  - Case "ScanState_moveActiveToInactive".  apply IHst. assumption.
  - Case "ScanState_moveActiveToHandled".   apply IHst. assumption.
  - Case "ScanState_moveInactiveToActive".  apply IHst. assumption.
  - Case "ScanState_moveInactiveToHandled". apply IHst. assumption.
Defined.

Lemma ScanState_more_unhandledExtent `(st : ScanState sd)
  (H : length (unhandled sd) > 1) :
  intervalExtent (projT2 (getInterval sd
                  (safe_hd (unhandled sd) (gt_one_gt_zero _ H)))) <
  unhandledExtent sd.
Proof.
  pose proof st as Hi0.
  apply ScanState_unhandledExtent in Hi0.
  ScanState_cases (induction st) Case; simpl in *.
  - Case "ScanState_nil". inversion H.
  - Case "ScanState_newUnhandled".
    clear IHst.
    apply ScanState_unhandledExtent in st.
    rename st into Hi.
    cmp_reflexive.
    destruct unh eqn:Heqe. inversion H. inversion H2.
    inversion Hi; inversion H1. inversion H2.
    simpl in *.
    specialize (H3 f).
    assert (forall n m, m > 0 -> n < m + n).
      intros. omega. apply H4. clear H4.
    inversion H3; inversion H4.
      pose (Interval_extent_nonempty (projT2 (geti f))). omega.
    omega.
  - Case "ScanState_dropUnhandled".
    clear IHst.
    apply ScanState_unhandledExtent in st.
    rename st into Hi.
    destruct unh eqn:Heqe. inversion H.
    subst. simpl in *.
    destruct l. inversion H. inversion H1.
    inversion Hi0; inversion H0.
      inversion H1.
    specialize (H2 f).
    inversion H2. inversion H3. inversion H4.
    inversion H3. omega.
  - Case "ScanState_moveActiveToInactive".  apply IHst. assumption.
  - Case "ScanState_moveActiveToHandled".   apply IHst. assumption.
  - Case "ScanState_moveInactiveToActive".  apply IHst. assumption.
  - Case "ScanState_moveInactiveToHandled". apply IHst. assumption.
Defined.

Definition nextUnhandled `(st : ScanState sd)
  : option { sd' : ScanStateDesc &
             { st' : ScanState sd' &
               CurrentInterval st' & SSMorphSt sd sd' } }.
Proof.
  pose (ScanState_sole_unhandledExtent st).
  pose (ScanState_more_unhandledExtent st).

  destruct sd.
  destruct unhandled0.
    apply None.
  apply Some.

  assert { xe : nat & unhandledExtent0 =
                      intervalExtent (projT2 (getInterval0 i)) + xe } as Hxe.
    exists (unhandledExtent0 - intervalExtent (projT2 (getInterval0 i))).
    apply Minus.le_plus_minus. subst. simpl in *.
    apply Lt.le_lt_or_eq_iff.
    destruct unhandled0.
      right. apply e. auto.
    left. apply l. simpl. omega.

  assert (unhandledExtent0 > 0) as Hu.
    apply (@ScanState_unhandledExtent_nonzero
           {| nextInterval := nextInterval0
            ; unhandledExtent := unhandledExtent0
            ; unhandled := i :: unhandled0
            ; active := active0
            ; inactive := inactive0
            ; handled := handled0
            ; getInterval := getInterval0
            ; assignments := assignments0
            ; unhandled_sorted := unhandled_sorted0
            ; lists_are_unique := lists_are_unique0 |}); simpl.
      apply st.
    omega.

  destruct Hxe. subst.
  pose (ScanState_dropUnhandled
        nextInterval0
        x i unhandled0
        unhandled_sorted0
        active0
        inactive0
        handled0
        getInterval0
        assignments0
        lists_are_unique0 st).

  eexists.
  pose (intervalExtent (projT2 (getInterval0 i))).
  exists s.

  rapply Build_CurrentInterval.
    apply i.
    apply (projT2 (getInterval0 i)).

  (* Prove that a call to [nextUnhandled] must always reduce the unhandled
     extent. *)
  clear s.
  constructor.
    constructor; auto.
    simpl. unfold intervalExtent.
    unfold intervalStart, intervalEnd.
    remember (getInterval0 i) as v.
    destruct v. simpl. omega.

  (* jww (2014-09-19): How can I remove this duplication? *)
  simpl. unfold intervalExtent.
  unfold intervalStart, intervalEnd.
  remember (getInterval0 i) as v.
  destruct v. simpl.
  assert (ibeg x0 < iend x0)
    by (apply (interval_nonempty x0)).
  apply lt_minus in H. omega.
Defined.

Definition moveActiveToHandled `(st : ScanState sd) `(x : IntervalId sd)
  (H : In x (active sd))
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' }.
Proof.
  pose (ScanState_moveActiveToHandled sd x st H). eexists. apply s.
  destruct sd. simpl.
  rapply Build_SSMorph; auto.
  apply Le.le_n_Sn.
Defined.

Definition moveActiveToHandled' `(st : ScanState sd) `(x : IntervalId sd)
  (H : In x (active sd))
  : { sd' : ScanStateDesc & ScanState sd' }.
Proof.
  pose (ScanState_moveActiveToHandled sd x st H). eexists. apply s.
Defined.

Definition moveActiveToInactive `(st : ScanState sd) `(x : IntervalId sd)
  (H : In x (active sd))
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' }.
Proof.
  pose (ScanState_moveActiveToInactive sd x st H). eexists. apply s.
  destruct sd. simpl.
  rapply Build_SSMorph; auto.
Defined.

Definition moveInactiveToActive `(st : ScanState sd) `(x : IntervalId sd)
  (H : In x (inactive sd))
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' }.
Proof.
  pose (ScanState_moveInactiveToActive sd x st H). eexists. apply s.
  destruct sd. simpl.
  rapply Build_SSMorph; auto.
Defined.

Definition moveInactiveToHandled `(st : ScanState sd) `(x : IntervalId sd)
  (H : In x (inactive sd))
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' }.
Proof.
  pose (ScanState_moveInactiveToHandled sd x st H). eexists. apply s.
  destruct sd. simpl.
  rapply Build_SSMorph; auto.
  apply Le.le_n_Sn.
Defined.

(* We need to know that [x] is not already a member of the [ScanState].  We
   know it was removed from the [ScanState] by [nextUnhandled], but it may
   have been split and the other parts added back to the unhandled list, so we
   need to know that it's not going to recur. *)
Definition addToActive `(st : ScanState sd) `(result : CurrentInterval st)
  (reg : PhysReg) : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' }.
Proof.
Admitted.
(*
  destruct st.
  destruct result.
  eexists {| nextInterval := nextInterval0
           ; unhandled    := unhandled0
           ; active       := currentIntervalId0 :: active0
           ; inactive     := inactive0
           ; handled      := handled0
           ; getInterval  := getInterval0
           ; assignments  := fun i =>
               if cmp_eq_dec i currentIntervalId0
               then Some reg
               else assignments0 i
           |}.
  rapply Build_SSMorph; simpl; auto.
  Grab Existential Variables.
  apply NoDup_swap.
  rewrite <- app_comm_cons.
  apply NoDup_swap_cons.
  apply NoDup_cons; assumption.
Defined.
*)

(** ** Main functions *)

Definition getRegisterIndex `(st : ScanState sd) (k : IntervalId sd -> nat)
  (z : PhysReg -> option nat) (is : list (IntervalId sd))
  : PhysReg -> option nat :=
  fold_right
    (fun x f => fun r =>
       match assignments sd x with
       | None => f r
       | Some a => if cmp_eq_dec a r then Some (k x) else f r
       end) z is.

Definition nextIntersectionWith `(st : ScanState sd)
  `(x : Interval xd) (yid : IntervalId sd) : nat.
Proof.
Admitted.

Function findRegister (freeUntilPos : PhysReg -> option nat) (reg : PhysReg)
  {measure fin_to_nat reg} : (PhysReg * option nat)%type :=
  match freeUntilPos reg with
  | None => (reg, None)
  | Some pos =>
      match pred_fin reg with
      | None => (reg, Some pos)
      | Some nreg =>
          match findRegister freeUntilPos nreg with
          | (reg', None) => (reg', None)
          | (reg', Some pos') =>
              if pos <? pos'
              then (reg', Some pos')
              else (reg,  Some pos)
          end
      end
  end.
Proof. intros. apply pred_fin_lt. assumption. Qed.

(** If [tryAllocateFreeReg] fails to allocate a register, the [ScanState] is
    left unchanged.  If it succeeds, or is forced to split [current], then a
    register will have been assigned. *)
Definition tryAllocateFreeReg `(st : ScanState sd) `(i : CurrentInterval st)
  : option (PhysReg *
            { sd' : ScanStateDesc &
              { st' : ScanState sd' &
                      CurrentInterval st' & SSMorph sd sd' } }) :=
  (* The first part of this algorithm has been modified to be more functional:
     instead of mutating an array called [freeUntilPos] and finding the
     register with the highest value, we use a function produced by a fold,
     and iterate over the register set. *)
  let currentId := currentIntervalId i in
  let cd        := currentDesc i in
  let current   := currentInterval i in

  (* set freeUntilPos of all physical registers to maxInt
     for each interval it in active do
       freeUntilPos[it.reg] = 0 *)
  let freeUntilPos' :=
        getRegisterIndex st (const 0) (const None) (active sd) in

  (* for each interval it in inactive intersecting with current do
       freeUntilPos[it.reg] = next intersection of it with current *)
  let intersectingIntervals :=
        filter (fun x => anyRangeIntersects
                           (rds cd) (rds (projT1 (getInterval sd x))))
               (inactive sd) in
  let freeUntilPos :=
        getRegisterIndex st (nextIntersectionWith st current) freeUntilPos'
                         intersectingIntervals in

  (* reg = register with highest freeUntilPos *)
  let lastReg     := ultimate_from_nat maxReg registers_exist in
  let (reg, mres) := findRegister freeUntilPos lastReg in
  let result      := existT _ sd (existT2 _ _ st i (newSSMorph sd)) in
  let useReg      := (reg, result) in

  (* [mres] indicates the highest use position of the indicated register,
     which is the furthest available. *)
  match mres with
  | None => Some useReg
  | Some n =>
      (* if freeUntilPos[reg] = 0 then
           // no register available without spilling
           allocation failed
         else if current ends before freeUntilPos[reg] then
           // register available for the whole interval
           current.reg = reg
         else
           // register available for the first part of the interval
           current.reg = reg
           split current before freeUntilPos[reg] *)
      if beq_nat n 0
      then None
      else if ltb (intervalEnd current) n
           then Some useReg
           else None            (* jww (2014-09-12): NYI *)
  end.

(** If [allocateBlockedReg] fails, it's possible no register was assigned and
    that the only outcome was to split one or more intervals.  This is why the
    type differs from [tryAllocateFreeReg], since in all cases the final state
    is changed. *)
Definition allocateBlockedReg `(st : ScanState sd) `(i : CurrentInterval st)
  : option PhysReg *
    { sd' : ScanStateDesc &
      { st' : ScanState sd' & CurrentInterval st' & SSMorph sd sd' } } :=
  (* set nextUsePos of all physical registers to maxInt *)

  (* for each interval it in active do
       nextUsePos[it.reg] = next use of it after start of current
     for each interval it in inactive intersecting with current do
       nextUsePos[it.reg] = next use of it after start of current *)

  (* reg = register with highest nextUsePos
     if first usage of current is after nextUsePos[reg] then
       // all other intervals are used before current, so it is best
       // to spill current itself
       assign spill slot to current
       split current before its first use position that requires a register
     else
       // spill intervals that currently block reg
       current.reg = reg
       split active interval for reg at position
       split any inactive interval for reg at the end of its lifetime hole *)

  (* // make sure that current does not intersect with
     // the fixed interval for reg
     if current intersects with the fixed interval for reg then
       split current before this intersection *)

  let result := existT _ sd (existT2 _ _ st i (newSSMorph sd)) in
  (None, result).

Definition activeIntervals `(st : ScanState sd)
  : list { i : IntervalId sd & In i (active sd) } :=
  let fix go l :=
      match l with
      | nil => nil
      | cons x xs =>
          existT _ x (in_eq x xs) :: map existT_in_cons (go xs)
      end in
  go (active sd).

(* Given a starting [ScanState] (at which point, [st = st0]), walk through the
   list of active intervals and mutate [st0] until it reflects the desired end
   state. *)
Fixpoint checkActiveIntervals `(st : ScanState sd) pos
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' } :=
  let fix go (sd : ScanStateDesc) (st : ScanState sd) ss is pos :=
    match is with
    | nil => ss
    | x :: xs =>
        (* // check for intervals in active that are handled or inactive
           for each interval it in active do
             if it ends before position then
               move it from active to handled
             else if it does not cover position then
               move it from active to inactive *)
        let i := projT2 (getInterval sd (projT1 x)) in
        let st1 := if intervalEnd i <? pos
                   then moveActiveToHandled st (projT1 x) (projT2 x)
                   else if negb (intervalCoversPos i pos)
                        then moveActiveToInactive st (projT1 x) (projT2 x)
                        else ss in
        go sd st st1 xs pos
    end in
  go sd st (existT2 _ _ sd st (newSSMorph sd)) (activeIntervals st) pos.

Definition inactiveIntervals `(st : ScanState sd)
  : list { i : IntervalId sd & In i (inactive sd) } :=
  let fix go l :=
      match l with
      | nil => nil
      | cons x xs =>
          existT _ x (in_eq x xs) :: map existT_in_cons (go xs)
      end in
  go (inactive sd).

Fixpoint checkInactiveIntervals `(st : ScanState sd) pos
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd sd' } :=
  let fix go (sd : ScanStateDesc) (st : ScanState sd) ss is pos :=
    match is with
    | nil => ss
    | x :: xs =>
        (* // check for intervals in inactive that are handled or active
           for each interval it in active do
             if it ends before position then
               move it from active to handled
             else if it covers position then
               move it from active to inactive *)
        let i := projT2 (getInterval sd (projT1 x)) in
        let st1 := if intervalEnd i <? pos
                   then moveInactiveToHandled st (projT1 x) (projT2 x)
                   else if intervalCoversPos i pos
                        then moveInactiveToActive st (projT1 x) (projT2 x)
                        else ss in
        go sd st st1 xs pos
    end in
  go sd st (existT2 _ _ sd st (newSSMorph sd)) (inactiveIntervals st) pos.

Definition handleInterval `(st0 : ScanState sd0) `(i : CurrentInterval st0)
  : { sd' : ScanStateDesc & ScanState sd' & SSMorph sd0 sd' } :=
  (* position = start position of current *)
  let currentId := currentIntervalId i in
  let position  := intervalStart (currentInterval i) in

  (* // check for intervals in active that are handled or inactive
     for each interval it in active do
       if it ends before position then
         move it from active to handled
       else if it does not cover position then
         move it from active to inactive *)
  let sp1  := checkActiveIntervals st0 position in
  let cid1 := transportId (next_interval_increases (projTT3 sp1)) currentId in

  (* // check for intervals in inactive that are handled or active
     for each interval it in inactive do
       if it ends before position then
         move it from inactive to handled
       else if it covers position then
         move it from inactive to active *)
  let sp2  := checkInactiveIntervals (projTT2 sp1) position in
  let cid2 := transportId (next_interval_increases (projTT3 sp2)) cid1 in

  (* // find a register for current
     tryAllocateFreeReg
     if allocation failed then
       allocateBlockedReg *)
  let (mreg, result) :=
      match tryAllocateFreeReg st0 i with
      | Some (reg, result) => (Some reg, result)
      | None => allocateBlockedReg st0 i
      end in

  (* if current has a register assigned then
       add current to active *)
  match result with
  | existT sd3 (existT2 st3 current' ss3) =>
      match mreg with
      | Some reg =>
          let (sd4,st4,ss4) := addToActive st3 current' reg in
          existT2 _ _ sd4 st4 (transitivity ss3 ss4)
      | None => existT2 _ _ sd3 st3 ss3
      end
  end.

Function linearScan (sd : ScanStateDesc) (st : ScanState sd)
  {measure unhandledExtent sd} : { sd' : ScanStateDesc & ScanState sd' } :=
  (* while unhandled /= { } do
       current = pick and remove first interval from unhandled
       HANDLE_INTERVAL (current) *)
  match nextUnhandled st with
  | None => existT _ sd st
  | Some (existT sd1 (existT2 st1 i smorph1)) =>
    match handleInterval st1 i with
    | existT2 sd2 st2 smorph2 => linearScan sd2 st2
    end
  end.
Proof.
  (* We must prove that after every call to handleInterval, the total extent
     of the remaining unhandled intervals is less than it was before. *)
  intros.
  apply SSMorphSt_proj_unhandledExtent.
  apply compose_SSMorph_with_SSMorphSt with (sd2 := sd1); assumption.
Defined.

(****************************************************************************)

(** * Program graphs *)

(** Given a node graph of our low-level intermediate representation, where
    instructions are associated with virtual registers, compute the linear
    mapping to intervals. *)

Class Graph (a : Set) := {}.

Definition determineIntervals (g : Graph VirtReg)
  : { sd : ScanStateDesc & ScanState sd }.
Admitted.

Definition allocateRegisters (g : Graph VirtReg)
  : { sd : ScanStateDesc & ScanState sd } :=
  let (sd,st) := determineIntervals g in linearScan sd st.

End Allocator.
